.npn_bjt_common_emitter.vcc in 0 DC [12]
.Rc in vcc out [4.7k]
.Re in vcc 0 [1k]

.basedivider.Rb1 in vcc base [100k]
.Rb2 in base 0 [20k]

.Q1 in base 12 NPN1
.NPN1 NPN
.OP
.END

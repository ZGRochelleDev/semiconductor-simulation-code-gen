[NETLIST]
V1 in 0
R1 in n1 1k
C1 n1 0 100n
R2 n1 out 1k
C2 out 0 0
.ac dec 100Hz 1MHz
.print ac V(out)

.END

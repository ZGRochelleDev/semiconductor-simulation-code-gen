*MOS1
vdd in 0 DC 1
RD in out 1k 
NMOS1 in out in 0 0 0 1
.vin in 0 DC 0
.dc vin 0 5 0.1
.print dc V(out)
.end

COMPONENTS
    V1 DC 1.2V
    R1 220 ohms
    ZD5V6 5.6V
    RLOAD 1K ohms
END COMPONENTS

INITIAL CONDITIONS
    V1 = 1.2V, R1 = 220 ohm, ZD5V6 = 5.6V, RLOAD = 1K ohm
END INITIAL CONDITIONS

ANALYSIS
    .OP
    .AC 1MHz
    .DC 1kHz
    .TRAN 1s
    .PRINT VOUT
    .MEAS VOUT
.END

**divider_op**
I1 in 0 DC
R1 in out
.end

.zener_regulator
V1 in 12
R1 in out
.DZ out 0 5.6
.Rload out 0 1
.op
.print Vout
.end

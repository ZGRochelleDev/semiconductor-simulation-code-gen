M1: NMOS1(0 0 0 0)
M2: NMOS1(1 1 1 1)

Rref: 10K(0 0 1 0)
RL: 10K(-1 -1 1 0)

.END

*. op
V1 in 1
E1 out 0 in out 10
.R load 10k
.end

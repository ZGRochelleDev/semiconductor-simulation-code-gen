* npn_bjt_common_emitter
vcc in 0 DC 12
Rc in out 4.7k
Re in emit 1k
.Rb1 in base 100k 100k+20k
.Rb2 in base 20k
.Q1 in emit base 0 NPN1
.op
.print op V(out), V(base)
.end

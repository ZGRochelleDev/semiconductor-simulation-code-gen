V(0)
I1 = 2mA
R1 = 1k
.END

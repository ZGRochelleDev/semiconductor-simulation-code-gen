V1 DC 1V
E1 OUT 0 IN 0 10
RLOAD 10K
.END

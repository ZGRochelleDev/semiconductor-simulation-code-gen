plaintext
divider_op
V1 in -1000000 0 5
R1 out 10000 1
C1 out 10e-9 0
.end

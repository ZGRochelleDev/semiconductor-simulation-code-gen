plaintext
divider_op
V1 in -1000000 0 5
R1 -1000 0
C1 0 10e-9
.end
